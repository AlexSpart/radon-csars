
import <execution_loop.cdl>;
functions = {f1, f2, f3, f4};
fs = 4;

f1.calls = {f2, f3};
f2.calls = {}; 
f3.calls = {f4};
f4.calls = {f1};

@show fn[1];
@show fn[2];
@show fn[3];
@show fn[4];